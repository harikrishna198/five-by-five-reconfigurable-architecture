----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/18/2023 09:54:41 AM
-- Design Name: 
-- Module Name: TestBench - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use std.env.finish;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TestBench is
--  Port ( );
end TestBench;

architecture Behavioral of TestBench is
Signal A1,A2,A3,A4,A5,B1,B2,B3,B4,B5:  std_logic_vector(3 downto 0);
Signal SEL11,SEL12,SEL13,SEL14,SEL15,
SEL21,SEL22, SEL23, SEL24,SEL25,
SEL31, SEL32, SEL33, SEL34, SEL35,
SEL41, sel42, sel43, sel44, SEL45,
SEL51,sel52, sel53, sel54, SEL55:  std_logic_vector(4 downto 0);
Signal t11, t12, t19, t110,
 t21, t22, t29, t210,
 t31, t32,t33, t34,  t37, t38,t39, t310,
 t41, t42,t43, t44, t45, t46, t47, t48, t49, t410:  std_logic;
Signal f13, f14,f15, f16,f17, f18,
f23, f24,f25, f26,f27, f28,
 f35,f36:  std_logic_vector(1 downto 0);
Signal  z1,z2,z3,z4,z5 :  std_logic_vector(3 downto 0 );
begin
dut: entity work.Top_Box(str)
port map(A1 => A1,A2 => A2,A3 => A3,A4 => A4,A5 => A5,B1 =>B1,B2 =>B2,B3 =>B3,B4 =>B4,B5 =>B5,
SEL11 => SEL11,SEL12 => SEL12,SEL13 => SEL13,SEL14 => SEL14,SEL15 => SEL15,
SEL21 => SEL21,SEL22 => SEL22, SEL23 => SEL23, SEL24 => SEL24,SEL25 => SEL25,
SEL31 => SEL31, SEL32 => SEL32, SEL33 => SEL33, SEL34 => SEL34, SEL35 => SEL35,
SEL41=> SEL41, sel42 => SEL42, sel43 => SEL43, sel44 => SEL44, SEL45 => SEL45,
SEL51 => SEL51,sel52 => SEL52, sel53 => SEL53, sel54 => SEL54, SEL55 => SEL55,
t11 =>t11 , t12 =>t12, t19 =>t19, t110 =>t110,
t21 =>t21, t22 =>t22, t29 =>t29, t210 =>t210,
 t31 =>t31, t32 =>t32,t33 =>t33, t34 =>t34,  t37 =>t37, t38 =>t38,t39 =>t39, t310 =>t310,
 t41 =>t41, t42 =>t42,t43 =>t43, t44 =>t44, t45 =>t45, t46 =>t46, t47 =>t47, t48 =>t48, t49 =>t49, t410 =>t410,
f13 =>f13, f14 =>f14,f15 =>f15, f16 =>f16,f17 =>f17, f18 =>f18,
f23 =>f23, f24 =>f24,f25 =>f25, f26 =>f26,f27 =>f27, f28 =>f28,
 f35 =>f35,f36=>f36,
z1 =>z1,z2 =>z2,z3 =>z3,z4 =>z4,z5 =>z5);

stim:process
begin
A1 <= "1001";A2 <= "0100";A3 <= "0010";A4 <= "1111";A5 <= "0001";B1 <="0110";B2 <="0011";B3 <="0111";B4 <="1101";B5 <="0001";
SEL11 <="00000";SEL12 <= "00010";SEL13 <= "00000";SEL14 <="00001";SEL15 <= "00010";
SEL21 <= "10011";SEL22 <="00001"; SEL23 <= "00000"; SEL24 <= "00001";SEL25 <="10001";
SEL31 <="10011"; SEL32 <="00011"; SEL33 <="00100"; SEL34 <="00101"; SEL35 <="10011";
SEL41<="10011"; sel42 <="00110"; sel43 <="10011"; sel44 <="01000"; SEL45 <="10011";
SEL51 <="10011";sel52 <="10001"; sel53 <="10011"; sel54 <="10010"; SEL55 <="10011";
t11 <='1'; t12 <='1';f13 <="01"; f14 <="10";f15 <="10"; f16 <="11";f17 <="00"; f18 <="10"; t19 <='1'; t110 <='0';
t21 <='1'; t22 <='0';f23 <="10"; f24 <="11";f25 <="10"; f26 <="10";f27 <="00"; f28 <="10"; t29 <='0'; t210 <='0';
t31 <='1'; t32 <='0';t33 <='1'; t34 <='1';f35<="10";f36<="10"; t37 <='0'; t38 <='0';t39 <='0'; t310 <='0';
 t41 <='1'; t42 <='0';t43 <='1'; t44 <='0'; t45 <='0'; t46 <='0'; t47 <='1'; t48 <='0'; t49 <='0'; t410 <='0';

 wait FOR 100NS;

A1 <= "1101";A2 <= "0010";A3 <= "0000";A4 <= "0001";A5 <= "0010";B1 <="0110";B2 <="0011";B3 <="0000";B4 <="0001";B5 <="0010";
SEL11 <="00001";SEL12 <= "00010";SEL13 <= "10011";SEL14 <="00000";SEL15 <= "00010";
SEL21 <= "10001";SEL22 <="00000"; SEL23 <= "00001"; SEL24 <= "00000";SEL25 <="10001";
SEL31 <="10011"; SEL32 <="01100"; SEL33 <="10000"; SEL34 <="10001"; SEL35 <="10011";
SEL41<="10011"; sel42 <="01001"; sel43 <="01011"; sel44 <="10011"; SEL45 <="10011";
SEL51 <="10011";sel52 <="10001"; sel53 <="10001"; sel54 <="10011"; SEL55 <="10011";
t11 <='1'; t12 <='0';f13 <="01"; f14 <="11";f15 <="00"; f16 <="11";f17 <="00"; f18 <="10"; t19 <='0'; t110 <='0';
t21 <='1'; t22 <='0';f23 <="00"; f24 <="11";f25 <="01"; f26 <="11";f27 <="01"; f28 <="00"; t29 <='0'; t210 <='0';
t31 <='1'; t32 <='0';t33 <='1'; t34 <='1';f35<="01";f36<="10"; t37 <='0'; t38 <='0';t39 <='0'; t310 <='0';
t41 <='1'; t42 <='1';t43 <='1'; t44 <='0'; t45 <='0'; t46 <='0'; t47 <='1'; t48 <='0'; t49 <='0'; t410 <='0';

 wait FOR 100NS;


A1 <= "1000";A2 <= "1110";A3 <= "0000";A4 <= "0001";A5 <= "0011";B1 <="0101";B2 <="1000";B3 <="0000";B4 <="0100";B5 <="0010";
SEL11 <="00000";SEL12 <= "00001";SEL13 <= "10011";SEL14 <="00010";SEL15 <= "00010";
SEL21 <= "10011";SEL22 <="00001"; SEL23 <= "00000"; SEL24 <= "00001";SEL25 <="10001";
SEL31 <="10011"; SEL32 <="10011"; SEL33 <="01000"; SEL34 <="00101"; SEL35 <="10011";
SEL41<="10011"; sel42 <="10011"; sel43 <="10001"; sel44 <="10001"; SEL45 <="10011";
SEL51 <="10011";sel52 <="10011"; sel53 <="10001"; sel54 <="10001"; SEL55 <="10011";
t11 <='1'; t12 <='0';f13 <="01"; f14 <="01";f15 <="00"; f16 <="11";f17 <="00"; f18 <="10"; t19 <='0'; t110 <='0';
t21 <='1'; t22 <='0';f23 <="01"; f24 <="01";f25 <="00"; f26 <="11";f27 <="01"; f28 <="01"; t29 <='0'; t210 <='0';
t31 <='1'; t32 <='0';t33 <='1'; t34 <='0';f35<="10";f36<="01"; t37 <='1'; t38 <='0';t39 <='0'; t310 <='0';
t41 <='1'; t42 <='1';t43 <='1'; t44 <='0'; t45 <='1'; t46 <='0'; t47 <='1'; t48 <='0'; t49 <='0'; t410 <='0';

 wait FOR 100NS;


A1 <= "0100";A2 <= "0011";A3 <= "0000";A4 <= "1111";A5 <= "0010";B1 <="0010";B2 <="0100";B3 <="0000";B4 <="1010";B5 <="0010";
SEL11 <="00010";SEL12 <= "00000";SEL13 <= "10011";SEL14 <="00001";SEL15 <= "00010";
SEL21 <= "10011";SEL22 <="00000"; SEL23 <= "00000"; SEL24 <= "00001";SEL25 <="10011";
SEL31 <="10011"; SEL32 <="01111"; SEL33 <="01101"; SEL34 <="01110"; SEL35 <="10011";
SEL41<="10011"; sel42 <="00110"; sel43 <="00111"; sel44 <="10011"; SEL45 <="10011";
SEL51 <="10011";sel52 <="01010"; sel53 <="10011"; sel54 <="10011"; SEL55 <="10011";
t11 <='1'; t12 <='0';f13 <="01"; f14 <="11";f15 <="01"; f16 <="11";f17 <="10"; f18 <="10"; t19 <='0'; t110 <='0';
t21 <='1'; t22 <='0';f23 <="10"; f24 <="10";f25 <="01"; f26 <="10";f27 <="01"; f28 <="01"; t29 <='0'; t210 <='0';
t31 <='1'; t32 <='0';t33 <='1'; t34 <='1';f35<="10";f36<="10"; t37 <='1'; t38 <='0';t39 <='0'; t310 <='0';
t41 <='1'; t42 <='1';t43 <='1'; t44 <='1'; t45 <='1'; t46 <='0'; t47 <='1'; t48 <='0'; t49 <='0'; t410 <='0';

 wait FOR 100NS;

 finish;
end process;
end Behavioral;
